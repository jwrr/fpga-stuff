module waves();
  initial begin
    $dumpfile(`VCD_OUT);
    $dumpvars(0, iceZ0mb1e);
  end
endmodule

